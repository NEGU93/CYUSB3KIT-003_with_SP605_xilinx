----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:40:48 12/11/2018 
-- Design Name: 
-- Module Name:    counter - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity counter is
    Port ( CLOCK : in  STD_LOGIC;
           DIRECTION : in  STD_LOGIC;
           COUNT_OUT : out  STD_LOGIC_VECTOR (3 downto 0)
			  );
end counter;

architecture Behavioral of counter is
signal count_int : std_logic_vector(3 downto 0) := "0000";
signal delayed_int : std_logic_vector(23 downto 0) := "000000000000000000000000";
begin
process(CLOCK)
begin
	if CLOCK='1' and CLOCK'event then
		if delayed_int = "000000000000000000000000" then
			if DIRECTION='1' then
				count_int <= count_int + 1;
			else
				count_int <= count_int - 1;
			end if;
		end if;
		delayed_int <= delayed_int + 1;
	end if;
end process;

COUNT_OUT <= count_int;
end Behavioral;
